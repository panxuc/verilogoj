module One(
    output out
);
    assign out = 1;
endmodule