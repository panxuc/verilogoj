module Zero(
    output out
);
    assign out = 0;
endmodule